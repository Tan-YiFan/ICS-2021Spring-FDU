`ifndef __PKG_SVH
`define __PKG_SVH

`include "common.sv"
`include "decode_pkg.sv"
`include "execute_pkg.sv"
`include "fetch_pkg.sv"
`include "forward_pkg.sv"
`include "memory_pkg.sv"
`include "writeback_pkg.sv"

`endif
