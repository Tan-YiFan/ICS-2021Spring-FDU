`include "mycpu/interface.svh"
module divider (
        
);
endmodule
